`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:23:48 05/17/2018 
// Design Name: 
// Module Name:    bancRegistres 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bancRegistres(
    input [15:0] A_no,
    input [15:0] B_no,
    input [15:0] W_no,
    input [15:0] Data,
    input W_flag,
    output [15:0] AS,
    output [15:0] BS
    );


endmodule
